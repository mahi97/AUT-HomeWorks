--------------------------------------------------------------------------------
-- Author:        Mohammad Mahdi Rahimi (mohammadmahdi76@gmail.com)
--
-- Create Date:   20-04-2017
-- Module Name:   ALU.vhd
--------------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
entity InstructionRegister is
  port (
	clock
  ) ;
end entity ; -- InstructionRegister

architecture arch of InstructionRegister is



begin



end architecture ; -- arch