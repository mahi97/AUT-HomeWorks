--------------------------------------------------------------------------------
-- Author:        Mohammad Mahdi Rahimi (mohammadmahdi76@gmail.com)
--
-- Create Date:   20-04-2017
-- Module Name:   ALU.vhd
--------------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
entity RegisterFile is
  port (
	clock
  ) ;
end entity ; -- RegisterFile

architecture behav of RegisterFile is



begin



end architecture ; -- behav