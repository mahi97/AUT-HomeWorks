--------------------------------------------------------------------------------
-- Author:        Mohammad Mahdi Rahimi (mohammadmahdi76@gmail.com)
--
-- Create Date:   20-04-2017
-- Module Name:   SAYEH.vhd
--------------------------------------------------------------------------------
library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
entity SAYEH is
  port (
	clock
  ) ;
end entity ; -- SAYEH

architecture behav of SAYEH is



begin



end architecture ; -- behav